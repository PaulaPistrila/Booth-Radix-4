library verilog;
use verilog.vl_types.all;
entity \_reg_file_tb\ is
end \_reg_file_tb\;
