library verilog;
use verilog.vl_types.all;
entity \_testbench\ is
end \_testbench\;
