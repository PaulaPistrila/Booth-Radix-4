library verilog;
use verilog.vl_types.all;
entity parallel_adder_tb is
end parallel_adder_tb;
